library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity cpu is
    Port(clk, rst, slct, start : in std_logic);
end cpu;

architecture Behavioral of cpu is

begin


end Behavioral;
