LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY cpu IS
    PORT (clk, rst, slct, start : IN STD_LOGIC);
END cpu;

ARCHITECTURE Behavioral OF cpu IS

BEGIN
END Behavioral;